.MODEL BC550_Cordell npn IS=45f BF=689 VAF=162 IKF=0.09 ISE=4600f NE=2 NF=0.9965 RB=167 RC=1 RE=0.04 CJE=18.7p MJE=0.35 VJE=0.75 CJC=6.2p MJC=0.25 VJC=0.4 FC=0.5 TF=595p XTF=10 VTF=10 ITF=1 TR=10n BR=12.2 IKR=0.34 EG=1.2 XTB=1.65 XTI=3 NC=0.996 NR=1.0 VAR=120 IRB=7e-5 RBM=1.1 XCJC=0.6 ISC=5f mfg=CA030111

.MODEL BC550B NPN(IS=1.8E-14 ISE=5.0E-14 ISC=1.72E-13 XTI=3 BF=400 BR=35.5 IKF=0.14 IKR=0.03 XTB=1.5 VAF=80 VAR=12.5 VJE=0.58 VJC=0.54 RE=0.6 RC=0.25 RB=0.56 CJE=13p CJC=4p XCJC=0.75 FC=0.5 NF=0.9955 NR=1.005 NE=1.46 NC=1.27 MJE=0.33 MJC=0.33 TF=0.64n TR=50.72n EG=1.11 VCEO=50 ICRATING=100M MFG=ZETEX)

.model BC550C NPN(Is=7.049f Xti=3 Eg=1.11 Vaf=23.89 Bf=493.2 Ise=99.2f Ne=1.829 Ikf=.1542 Nk=.6339 Xtb=1.5 Br=2.886 Isc=7.371p Nc=1.508 Ikr=5.426 Rc=1.175 Cjc=5.5p Mjc=.3132 Vjc=.4924 Fc=.5 Cje=11.5p Mje=.6558 Vje=.5 Tr=10n Tf=420.3p Itf=1.374 Xtf=39.42 Vtf=10 Vceo=30 Icrating=100m mfg=Philips)

.MODEL BC560A PNP(IS=1.149E-14 ISE=5E-14 ISC=1.43E-14 XTI=3 BF=330 BR=13 IKF=0.1 IKR=0.012 XTB=1.5 VAF=84.56 VAR=8.15 VJE=0.65 VJC=0.565 RE=0.4 RC=0.95 RB=0.2 CJE=16p CJC=10.5p XCJC=0.75 FC=0.5 NF=0.9872 NR=0.996 NE=1.4 NC=1.1 MJE=0.415 MJC=0.415 TF=0.493n TR=73.55n EG=1.11 VCEO=45V ICRATING=100M MFG=ZETEX)

.model BC560B PNP(Is=1.02f Xti=3 Eg=1.11 Vaf=51.26 Bf=289.6 Ise=9.846f Ne=1.845 Ikf=.1026 Nk=.5413 Xtb=1.5 Br=6.124 Isc=1.113f Nc=1.97 Ikr=.2035 Rc=1.078 Cjc=9.81p Mjc=.332 Vjc=.4865 Fc=.5 Cje=30p Mje=.3333 Vje=.5 Tr=10n Tf=612.4p Itf=1.287 Xtf=25.55 Vtf=10 Vceo=30 Icrating=100m mfg=Philips)

.model BC560C PNP(Is=1.02f Xti=3 Eg=1.11 Vaf=34.62 Bf=401.6 Ise=38.26p Ne=5.635 Ikf=74.73m Nk=.512 Xtb=1.5 Br=9.011 Isc=1.517f Nc=1.831 Ikr=.1469 Rc=1.151 Cjc=9.81p Mjc=.332 Vjc=.4865 Fc=.5 Cje=30p Mje=.3333 Vje=.5 Tr=10n Tf=524p Itf=.9847 Xtf=17.71 Vtf=10 Vceo=30 Icrating=100m mfg=Philips)

.MODEL BC560_Cordell pnp IS=60f BF=900 VAF=160 IKF=0.10 ISE=70f NE=1.42 NF=1 RB=170 RC=1.0 RE=0.05 CJE=19p MJE=0.3 VJE=0.75 CJC=3.9p MJC=0.3 VJC=0.75 FC=0.5 TF=600p XTF=7 VTF=4 ITF=0.45 TR=10n BR=3 IKR=0 EG=1.1 XTB=1.5 XTI=3 NC=2 ISC=0 mfg=CA030211

.model 2N2222 NPN(IS=1E-14 VAF=100 BF=200 IKF=0.3 XTB=1.5 BR=3 CJC=8E-12 CJE=25E-12 TR=100E-9 TF=400E-12 ITF=1 VTF=2 XTF=3 RB=10 RC=.3 RE=.2 Vceo=30 Icrating=800m mfg=Philips)
